library verilog;
use verilog.vl_types.all;
entity adderTB is
end adderTB;
