library verilog;
use verilog.vl_types.all;
entity adderDoubleTB is
end adderDoubleTB;
