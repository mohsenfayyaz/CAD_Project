library verilog;
use verilog.vl_types.all;
entity single_divider_TB is
end single_divider_TB;
