library verilog;
use verilog.vl_types.all;
entity Main_TB_2_corner_case is
end Main_TB_2_corner_case;
