library verilog;
use verilog.vl_types.all;
entity double_divider_TB is
end double_divider_TB;
