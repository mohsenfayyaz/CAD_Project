library verilog;
use verilog.vl_types.all;
entity double_adder_TB is
end double_adder_TB;
