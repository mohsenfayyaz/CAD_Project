library verilog;
use verilog.vl_types.all;
entity sqrtTB is
end sqrtTB;
