library verilog;
use verilog.vl_types.all;
entity multiplier_TB is
end multiplier_TB;
