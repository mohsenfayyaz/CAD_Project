library verilog;
use verilog.vl_types.all;
entity double_multiplier_TB is
end double_multiplier_TB;
