library verilog;
use verilog.vl_types.all;
entity multiplierTB is
end multiplierTB;
