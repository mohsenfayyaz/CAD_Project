library verilog;
use verilog.vl_types.all;
entity single_sqrt_TB is
end single_sqrt_TB;
