library verilog;
use verilog.vl_types.all;
entity Main_TB is
end Main_TB;
