library verilog;
use verilog.vl_types.all;
entity Main_TB_2 is
end Main_TB_2;
