library verilog;
use verilog.vl_types.all;
entity dividerTB is
end dividerTB;
