library verilog;
use verilog.vl_types.all;
entity double_sqrt_TB is
end double_sqrt_TB;
